$display("%-15s%-10s%-10s%-10s%-10d%-10d%-10d%-10d%-10d%-15d%-10d%-10d%-10d",
{state_str},
{ty_str},
{pe_x_str},
{pe_y_str},
dut.sub_placer_{ty}_inst.pe_x{x}_y{y}.blk_id,
dut.sub_placer_{ty}_inst.pe_x{x}_y{y}.X,
dut.sub_placer_{ty}_inst.pe_x{x}_y{y}.Y,
dut.sub_placer_{ty}_inst.pe_x{x}_y{y}.sum_px,
dut.sub_placer_{ty}_inst.pe_x{x}_y{y}.sum_py,
dut.sub_placer_{ty}_inst.pe_x{x}_y{y}.temp_blk_id,
dut.sub_placer_{ty}_inst.pe_x{x}_y{y}.temp_coord[2*$clog2({B_t} + 1) - 1:$clog2({B_t} + 1)],
dut.sub_placer_{ty}_inst.pe_x{x}_y{y}.temp_coord[$clog2({B_t} + 1) - 1:0],
dut.sub_placer_{ty}_inst.pe_x{x}_y{y}.temp);