module dummy_benchmark(input wire i, output wire o);

    assign o = i;

endmodule